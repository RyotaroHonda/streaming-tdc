library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package defGateGen is

  constant kWidthTrgDelay : integer:= 8;
  constant kWidthTrgWidth : integer:= 16;

end package;